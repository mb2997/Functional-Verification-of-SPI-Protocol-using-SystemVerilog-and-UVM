`define HDR_LEN 16
`define ADD_LEN 14
`define DLY_LEN 4
`define DATA_LEN 32
`define CYCLE 10
`define NO_DATA_WIDTH 3